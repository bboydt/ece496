module top (
    input clk30
)

endmodule;
